module SR_FF (
    input S, R, clk, rst, Q,  
    output reg Qn             
);

always @(posedge clk or posedge rst) begin
	if (rst) begin
            Qn <= 1'b0;  
        end else begin
            if (S && R) begin
                Qn <= 1'bx;  
            end else if (S) begin
                Qn <= 1'b1;  
            end else if (R) begin
                Qn <= 1'b0;  
            end else begin
                Qn <= Q;  
            end
        end
end    
endmodule    
