`timescale 1ps/1ps
module SR_FF_tb ();    
reg S, R, clk, rst, Q;
wire Qn;

SR_FF dut (
    .S(S),
    .R(R),
    .clk(clk),
    .rst(rst),
    .Q(Q),
    .Qn(Qn)
);
initial begin
    clk = 0;
    forever #5 clk = ~clk;
end

initial begin
    $monitor("S = %b, R = %b, Q = %b", S, R, Q);
    rst = 1;
    #10 rst = 0;
    Q = 1;
    S = 0; R = 0; #10;
    S = 1; R = 0; #10;
    S = 0; R = 1; #10;
    S = 1; R = 1; #10;
    S = 0; R = 0; #10;
    $finish;
end

endmodule