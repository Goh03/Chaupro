module T_FF (
    input T,clk,
    

);
    
endmodule